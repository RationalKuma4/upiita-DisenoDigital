library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

entity Examen is Port
(
	clk   : IN  STD_LOGIC;
        reset : IN  STD_LOGIC;
        D0    : IN  STD_LOGIC_VECTOR(5 downto 0);
        D1    : IN  STD_LOGIC_VECTOR(5 downto 0);
        D2    : IN  STD_LOGIC_VECTOR(5 downto 0);
        D3    : IN  STD_LOGIC_VECTOR(5 downto 0);
        salida: OUT STD_LOGIC_VECTOR(7 downto 0);
        MUX   : OUT STD_LOGIC_VECTOR(3 downto 0)
);
end Examen;

architecture Arq_Examen of Examen is
	COMPONENT clk200Hz IS
        PORT (
            entrada: IN  STD_LOGIC;
            reset  : IN  STD_LOGIC;
            salida : OUT STD_LOGIC
        );
    END COMPONENT;
     
    COMPONENT siete_segmentos IS
        PORT (
            entrada: IN  STD_LOGIC_VECTOR(5 downto 0);
            salida : OUT STD_LOGIC_VECTOR(7 downto 0)
        );
    END COMPONENT;
     
    COMPONENT siete_segmentos_mux IS
        PORT (
            clk   : IN  STD_LOGIC;
            reset : IN  STD_LOGIC;
            D0    : IN  STD_LOGIC_VECTOR(5 downto 0);
            D1    : IN  STD_LOGIC_VECTOR(5 downto 0);
            D2    : IN  STD_LOGIC_VECTOR(5 downto 0);
            D3    : IN  STD_LOGIC_VECTOR(5 downto 0);
            salida: OUT STD_LOGIC_VECTOR(5 downto 0);
            MUX   : OUT STD_LOGIC_VECTOR(3 downto 0)
        );
    END COMPONENT;
     
    signal clk_out : STD_LOGIC := '0';
    signal digito  : STD_LOGIC_VECTOR(5 downto 0);
begin
	clk_i: clk200Hz PORT MAP(
        clk, reset, clk_out
    );
     
    mux_i: siete_segmentos_mux PORT MAP(
        clk_out, reset, "000000", "000001", "000010", "000011", digito, MUX
    );
     
    seg_i: siete_segmentos PORT MAP(
        digito, salida
    );
end Arq_Examen;

