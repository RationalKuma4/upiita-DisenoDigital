----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:14:29 10/23/2016 
-- Design Name: 
-- Module Name:    VhdlPrueba - Arq_VhdlPrueba 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity VhdlPrueba is
    Port ( a : in  STD_LOGIC;
           b : in  STD_LOGIC;
           y : inout  STD_LOGIC);
end VhdlPrueba;

architecture Arq_VhdlPrueba of VhdlPrueba is

begin


end Arq_VhdlPrueba;

